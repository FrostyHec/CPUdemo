`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/12/27 11:04:45
// Design Name: 
// Module Name: vga_disp
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module vga_disp(  
    input wire [31:0] digit, // input digit to show
    
    input wire vga_clk, // the clock of vga
    input wire rst, // reset
    input wire [9:0] x_pix, // x pixel position
    input wire [9:0] y_pix, // y pixel position
    output reg [11:0] pix_data // rgb of the pixel
);

parameter h_range = 10'd640; // 640
parameter v_range = 10'd480; // 480

// color
parameter   red = 12'hF80,
            orange = 12'hFC0,
            yellow = 12'hFFE,
            green = 12'h07E,
            cyan = 12'h07F,
            blue = 12'h01F,
            purple = 12'hF81,
            black = 12'h000,
            white = 12'hFFF,
            gray = 12'hD69;
            
reg [2047:0] char;

parameter x_begin = 10'd160, x_end = 10'd480;
parameter y_begin = 10'd208, y_end = 10'd272;
parameter char_wid = 10'd32;

parameter zero = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007E000001FF800003C1E0000700F0000E0070001E0038003C003C003C001C0078001E0078000E0070000E00F0000F00F0000F00F0000F00F0000701E0000781E0000781E0000781E0000781E0000781E0000781E0000781E0000781E0000781E0000781E0000781E0000781E0000781E0000780F0000700F0000F00F0000F00F0000F0070000E0078001E0078001E003C001C003C003C001E0038000E0070000700F00003C1E00001FF8000007E000000000000000000000000000000000000000000000000000000000000000000000000000,
          one = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040000000C0000001C0000007C00001FFC00001FFC0000007C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000007E000000FF00001FFFF8001FFFF80000000000000000000000000000000000000000000000000000000000000000000000000,
          two = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF000003FFE0000F81F0001E0078003C003C0078001E0070001E0070000F00F0000F00F8000F00F8000F00FC000F00FC000F00FC000F0078001E0000001E0000001E0000003C0000003C00000078000000F0000000E0000001C0000003800000070000000E0000001C0000003800000070000000E0000001C0000003800000070000000E0003001C000300380003007800030070000600E0000E01C0001E01FFFFFE01FFFFFE01FFFFFE01FFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000,
          three = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FE000007FF80000E07C0001801E0003000F000300078007000780070007C0078003C0078003C0078003C0030003C0000003C0000003C0000007800000078000000F0000000E0000003C000000F800000FE000000FF80000007C0000000F0000000780000003C0000001C0000001E0000000E0000000F0000000F0000000F0038000F007C000F00FC000F00FC000F00FC001E00F8001E0078003C00780038003C0070001F01E00007FFC00001FE000000000000000000000000000000000000000000000000000000000000000000000000000,
          four = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000E0000000E0000001E0000003E0000003E0000007E000000FE000000DE0000019E0000039E0000031E0000071E0000061E00000C1E00001C1E0000181E0000301E0000701E0000601E0000C01E0001C01E0001801E0003001E0003001E0006001E000E001E000C001E0018001E0038001E003FFFFFFC3FFFFFFC00001E0000001E0000001E0000001E0000001E0000001E0000001E0000001E0000001E0000001E0000003F00000FFFF8000FFFF8000000000000000000000000000000000000000000000000000000000000000000000000,
          five = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FFFFE001FFFFE001FFFFE001FFFFC001800000018000000180000001800000018000000180000001800000018000000100000001000000030000000303F800031FFE00033FFF0003781F80036007C003C003C0038003E0038001E0000001E0000001F0000000F0000000F0000000F0000000F0000000F0000000F0038000F007C000F00FC000F00FC000E00FC001E00F8001E00F8001C0078003C00380078001C00F0000F01E00007FFC00000FE000000000000000000000000000000000000000000000000000000000000000000000000000,
          six = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FC000007FF00001E0780003803C0007003E000E003E001C003E0038003E0038001C00700000007000000070000000F0000000F0000000E0000000E0000000E03F8001E0FFF001E3FFF801E7C0FC01EF003E01EE001E01FC001F01F8000F01F0000F01F0000781E0000781E0000781E0000781E0000781E0000780E0000780F0000780F0000780F000070070000F0078000F003C000E003C001E001E001C000F00380007C0F00003FFE000007F000000000000000000000000000000000000000000000000000000000000000000000000000,
          seven = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFF007FFFFF007FFFFF007FFFFE007C000C0070000C006000180060001800C0003000C0003000C0006000000060000000C0000001C000000180000003800000038000000300000007000000070000000E0000000E0000001E0000001C0000003C0000003C00000038000000780000007800000078000000F8000000F8000000F8000000F8000000F8000001F8000001F8000001F8000001F8000001F8000001F8000001F8000001F8000000F0000000000000000000000000000000000000000000000000000000000000000000000000000,
          eight = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FF000007FFE0000F81F0001E0078003C003C0078001E0078001E00F0000F00F0000F00F0000F00F0000F00F0000F00F8000F00F8000E007C001E007E001C003F003C001FC078000FF0E00007FDC00001FF000003FF80000F1FE0001E07F0003C03F8007801FC0078007C00F0003E00F0003E01E0001F01E0001F01E0000F01E0000F01E0000F01E0000F01E0000F00F0000E00F0001E0078001C0078003C003E0078000F81F00007FFC00000FF000000000000000000000000000000000000000000000000000000000000000000000000000,
          nine = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001FE000007FF80000F03C0001E00E0003C0070007800380070003800F0001C00F0001C00E0001E01E0000E01E0000E01E0000E01E0000F01E0000F01E0000F01E0000F01E0000F01E0001F01F0001F00F0003F00F8006F00F800EF007C01CF003F07CF001FFF8F000FFE0F0003F81E0000001E0000001E0000001E0000001C0000003C0000003C0000003800380078007C0070007C00F0007C00E0007C01C0003C0380003E0F00001FFE000003F0000000000000000000000000000000000000000000000000000000000000000000000000000,
          ten = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003C0000003C0000003C0000007E0000007E0000006E0000006E000000CF000000CF000000C7000000C70000018780000187800001878000018380000303C0000303C0000303C0000301C0000601E0000601E0000601E0000600E0000E00E0000C00F0000C00F0000FFFF0001FFFF0001800780018007800180078003800780030003C0030003C0030003C0070003C0060001E0060001E0060001E00E0001E00E0001F01F0001F87FC00FFE7FC00FFE000000000000000000000000000000000000000000000000000000000000000000000000,
          eleven = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFF8003FFFFF0007C01F80078007C0078003E0078001E0078001F0078000F0078000F0078000F0078000F0078000F0078000F0078000E0078001E0078001E0078003C007800F0007801E0007FFF00007FFFC0007801F00078003C0078001E0078000F0078000700780007807800078078000380780003C0780003C0780003C0780003C0780003C0780003C0780003C0780007807800078078000F0078001F0078003E007C00FC07FFFFF007FFFF800000000000000000000000000000000000000000000000000000000000000000000000000,
          twelve = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FC10000FFFF0003C07F0007801F000E000F801C0007803C0003803800018078000180700000C0F00000C0E0000081E0000001E0000001E0000001E0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000001E0000001E0000001E0000081E00000C1E00000C0F0000080F000018078000100780003003C0006001E000C000F001C0007C0700001FFE000007F800000000000000000000000000000000000000000000000000000000000000000000000000,
          thirteen = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000007FFF80007FFFF0000FC07C0007801E0007800780078003C0078001C0078001E0078000F0078000F007800070078000780780007807800078078000380780003C0780003C0780003C0780003C0780003C0780003C0780003C0780003C0780003C0780003C0780003C0780003C0780003C0780003807800078078000780780007807800078078000F0078000F0078000E0078001E0078003C00780078007800F0007803E000FC0FC007FFFF0007FFF8000000000000000000000000000000000000000000000000000000000000000000000000000,
          fourteen = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFC03FFFFFE007E007E003C001E003C000F003C0007003C0003003C0003803C0001803C0000003C0000003C0000003C0060003C0060003C0060003C0060003C0060003C00E0003C01E0003FFFE0003FFFE0003C01E0003C00E0003C00E0003C0060003C0060003C0060003C0060003C0000003C0000003C0000003C0000003C0000003C0000003C0000C03C0000C03C0001803C0001803C0003803C0007803C000F007E003F03FFFFFF03FFFFFE0000000000000000000000000000000000000000000000000000000000000000000000000,
          fifteen = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000003FFFFFF03FFFFFF807E003F803C000F803C0003C03C0001C03C0000C03C0000E03C0000603C0000403C0000003C0000003C0000003C0000003C0030003C0030003C0030003C0030003C0070003C00F0003FFFF0003FFFF0003C00F0003C0070003C0070003C0030003C0030003C0030003C0030003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000003C0000007E000003FFC00003FFC0000000000000000000000000000000000000000000000000000000000000000000000000000,
          x = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000FFC3FF00FFC3FF001F0038000F0030000F0060000780E00003C0C00003C1800001E3800001E3000000F60000007E0000007C0000003C0000003C0000007E0000006F000000CF000001C78000018380000303C0000701E0000600E0000C00F0001C007800180078007C007E03FF03FF83FF03FF8000000000000000000000000000000000000000000000000000000000000000000000000;

reg [9:0] x_rel;
always@ (posedge vga_clk) begin
    x_rel = x_pix - x_begin;
    if (x_rel >= 0 && x_rel < char_wid * 1) begin
        char = zero;
    end
    else if (x_rel >= (char_wid * 1) && x_rel < (char_wid * 2)) begin
        char = x;
    end
    else if (x_rel >= (char_wid * 2) && x_rel < (char_wid * 3)) begin
        case(digit[31:28])
            4'b0000: char <= zero;
            4'b0001: char <= one;
            4'b0010: char <= two;
            4'b0011: char <= three;
            4'b0100: char <= four;
            4'b0101: char <= five;
            4'b0110: char <= six;
            4'b0111: char <= seven;
            4'b1000: char <= eight;
            4'b1001: char <= nine;
            4'b1010: char <= ten;
            4'b1011: char <= eleven;
            4'b1100: char <= twelve;
            4'b1101: char <= thirteen;
            4'b1110: char <= fourteen;
            4'b1111: char <= fifteen;
            default: char <= 2048'b0;
        endcase
    end
    else if (x_rel >= (char_wid * 3) && x_rel < (char_wid * 4)) begin
        case(digit[27:24])
            4'b0000: char <= zero;
            4'b0001: char <= one;
            4'b0010: char <= two;
            4'b0011: char <= three;
            4'b0100: char <= four;
            4'b0101: char <= five;
            4'b0110: char <= six;
            4'b0111: char <= seven;
            4'b1000: char <= eight;
            4'b1001: char <= nine;
            4'b1010: char <= ten;
            4'b1011: char <= eleven;
            4'b1100: char <= twelve;
            4'b1101: char <= thirteen;
            4'b1110: char <= fourteen;
            4'b1111: char <= fifteen;
            default: char <= 2048'b0;
        endcase
    end
    else if (x_rel >= (char_wid * 4) && x_rel < (char_wid * 5)) begin
        case(digit[23:20])
            4'b0000: char <= zero;
            4'b0001: char <= one;
            4'b0010: char <= two;
            4'b0011: char <= three;
            4'b0100: char <= four;
            4'b0101: char <= five;
            4'b0110: char <= six;
            4'b0111: char <= seven;
            4'b1000: char <= eight;
            4'b1001: char <= nine;
            4'b1010: char <= ten;
            4'b1011: char <= eleven;
            4'b1100: char <= twelve;
            4'b1101: char <= thirteen;
            4'b1110: char <= fourteen;
            4'b1111: char <= fifteen;
            default: char <= 2048'b0;
        endcase
    end
    else if (x_rel >= (char_wid * 5) && x_rel < (char_wid * 6)) begin
        case(digit[19:16])
            4'b0000: char <= zero;
            4'b0001: char <= one;
            4'b0010: char <= two;
            4'b0011: char <= three;
            4'b0100: char <= four;
            4'b0101: char <= five;
            4'b0110: char <= six;
            4'b0111: char <= seven;
            4'b1000: char <= eight;
            4'b1001: char <= nine;
            4'b1010: char <= ten;
            4'b1011: char <= eleven;
            4'b1100: char <= twelve;
            4'b1101: char <= thirteen;
            4'b1110: char <= fourteen;
            4'b1111: char <= fifteen;
            default: char <= 2048'b0;
        endcase
    end
    else if (x_rel >= (char_wid * 6) && x_rel < (char_wid * 7)) begin
        case(digit[15:12])
            4'b0000: char <= zero;
            4'b0001: char <= one;
            4'b0010: char <= two;
            4'b0011: char <= three;
            4'b0100: char <= four;
            4'b0101: char <= five;
            4'b0110: char <= six;
            4'b0111: char <= seven;
            4'b1000: char <= eight;
            4'b1001: char <= nine;
            4'b1010: char <= ten;
            4'b1011: char <= eleven;
            4'b1100: char <= twelve;
            4'b1101: char <= thirteen;
            4'b1110: char <= fourteen;
            4'b1111: char <= fifteen;
            default: char <= 2048'b0;
        endcase
    end   
    else if (x_rel >= (char_wid * 7) && x_rel < (char_wid * 8)) begin
        case(digit[11:8])
            4'b0000: char <= zero;
            4'b0001: char <= one;
            4'b0010: char <= two;
            4'b0011: char <= three;
            4'b0100: char <= four;
            4'b0101: char <= five;
            4'b0110: char <= six;
            4'b0111: char <= seven;
            4'b1000: char <= eight;
            4'b1001: char <= nine;
            4'b1010: char <= ten;
            4'b1011: char <= eleven;
            4'b1100: char <= twelve;
            4'b1101: char <= thirteen;
            4'b1110: char <= fourteen;
            4'b1111: char <= fifteen;
            default: char <= 2048'b0;
        endcase
    end
    else if (x_rel >= (char_wid * 8) && x_rel < (char_wid * 9)) begin
        case(digit[7:4])
            4'b0000: char <= zero;
            4'b0001: char <= one;
            4'b0010: char <= two;
            4'b0011: char <= three;
            4'b0100: char <= four;
            4'b0101: char <= five;
            4'b0110: char <= six;
            4'b0111: char <= seven;
            4'b1000: char <= eight;
            4'b1001: char <= nine;
            4'b1010: char <= ten;
            4'b1011: char <= eleven;
            4'b1100: char <= twelve;
            4'b1101: char <= thirteen;
            4'b1110: char <= fourteen;
            4'b1111: char <= fifteen;
            default: char <= 2048'b0;
        endcase
    end   
    else if (x_rel >= (char_wid * 9) && x_rel < (char_wid * 10)) begin
        case(digit[3:0])
            4'b0000: char <= zero;
            4'b0001: char <= one;
            4'b0010: char <= two;
            4'b0011: char <= three;
            4'b0100: char <= four;
            4'b0101: char <= five;
            4'b0110: char <= six;
            4'b0111: char <= seven;
            4'b1000: char <= eight;
            4'b1001: char <= nine;
            4'b1010: char <= ten;
            4'b1011: char <= eleven;
            4'b1100: char <= twelve;
            4'b1101: char <= thirteen;
            4'b1110: char <= fourteen;
            4'b1111: char <= fifteen;
            default: char <= 2048'b0;
        endcase
    end     
end

reg [9:0] x_pos;
reg [9:0] y_pos;

always@ (posedge vga_clk, negedge rst) begin
    if (rst == 1'b0) begin
        pix_data <= black;
    end
    else if(x_pix >= x_begin && x_pix <= x_end && y_pix >= y_begin && y_pix <= y_end) begin
        x_pos <= x_rel - x_rel / char_wid * char_wid;
        y_pos <= y_pix - y_begin;
        if(char[x_pos + y_pos * char_wid]) begin
            pix_data <= white;
        end
        else begin
            pix_data <= black;
        end
    end
    else begin
        pix_data <= black;
    end
end

endmodule
